BZh91AY&SYI��  �߀Px����߰?���P9�3dֵ��Q�M�j&j�� �4=@�9�&& &#4���d�#�����d�M y@h hb�2b`b0#L1&L0I�#	�0�<�Ѓ�  4�L(��*
�B��k%��ç�P�V��V�Z��M�5j�%�#�ƺ~
�t��?:����jTpy�"1���L#.�L(t�J�@c������([�׿È�(F���V��i[�i�#�5gq�����fP�h�!\��v��CN�����6�1��������#e$��z�Z�
�Y�+��?9g-`X5�[ޓK��ٿ�E����zss8��)�ӭ�u:jOE͗�WE�V����S0�Ѿ~�Z��%���	�vZӃ@kX~ ��DY��BF����/݆��1~��K�,w�h��`����}�X2���NZ1�{���T�e��ß��ޝ�\�E�P��b�&q�P��Gf�o"�=�vk�V�$� ��3Z��vl!��Li/C��+�9i���I:*�Weyj� `MN[�Dp�F�~�Es�eۆe����9\����y��w��9��Lŀ��+�����o�ט����E����5ݪUȪ(r��|b�L�*z�#�h���ys�	,�g�<��1���@q�E�Vlt?H)�+9�Ӌ��lV�s��ːDs���o6�R`�LI����#N(ϟ_�J/�&%f-:oW^��#�����7�	
 U��w#!��cZ���t�����)3#�\�K���fa@��;�]��BA$k׼