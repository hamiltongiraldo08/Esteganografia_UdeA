BZh91AY&SYD���  �߀Px����߰����P>��stk�p�S*6���6A�&���4i�hda��&��I��$��#A�@ 4   D�#Q5S���=P�  b �101��&$I�F�d�(i��@  ���YB{��AH)�[]��C`���(H�@nj�*�f��.��*{H�8�~�c�e�Bj�43��gV	�<��3PȨ֚F�L/��K< �,��*�E+h��˧pC&fG<�(�����=Ɂ��V������(�]Zf�w�
w��N�����ގ?�����l��+m��	Či?�ݔcw}0V����.Jl�����1632��Uo������fb�SD�5�Ug�T��ϴ_�?��}��2�,:Z7G�]�uUyy����]M\N�B� r��EA�\�)��#�1&+)+��\�E#��6�-܌V����v�X�9qWaES�ܜ则�R�Dg�O!�)Fã�~��H!���0��N�c��
_B?}�U�*\Q��m��Z�\�ޅ��g��DWj`chKRK�Ƹ|S�8�tך�Xi\���&��XW{T�)��K5'l�k�/ˈ���kc�4�wBf���Fyp�!g7����d�>sL��U6@ֹ*�$�ZI���&���l5��1$V�֬T���8�Eg��&�&`j�9]�Ԭ�!)`�T�3��D�U�4x�G��2f�*	
�
�AlfH�צ��myV�����Q\N�Ϭ�-*6	B��"x�h���p���R0�D��\��dz�(Ɉ^�61���F�w$S�	K�
�