BZh91AY&SYhI�  �߀Px����߰����P>wUq�:N��QL��zL�Se4=�i�h 2zC�4�H�ML����M��d� 2 4	M"bS�4��  � ѓ �`A��2`�DI2z�����<P4 h @V��!��J?�_�KC`�O�P�c@vڱ�cY��U�q�^�>�1���w34�d���o����h�β"/�DY�f6-n�)`�,x��;H�ѻ��;��^7`�a~;%���:a&	5m5�)�VR%�ѫH[޼5|��]��3&�331���5���?^i�B�\�l`F���/"�8���̠}��qU�̰���(�/�9y	�,y���i��&���\襳���h�5z���_1H�����q3��CQ~gd�9(+��-!D�̗��h�F&re*��Z�Q�"�N
^+P]�Ru�
��U��f�h�R��.��oT�X��A��^��>�@w}F+�;)X�OjĨ'=Q����J�/)�n�}�j�i�oB��3���8"�=� ʆ�.[�*t��G�M�H��#�PԻ&�[�M�]�+��3!(�k�k�O"�1�2���������&�D�x�!e �DFs���R�jzV32��R�� �'1L��_id(�7e� 6�Ó�AE��7;k���t9뉐8ǲ�|.��՜��%JrΒb&ATJk�.�7��-0������FPC�ْ5j��[e�qb�v�%�L�K�vV�G!;2  ����G�
��z����e���ř��e;�:B`Wy'�.�p� В?$